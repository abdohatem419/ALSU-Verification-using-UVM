package ALSU_main_sequence_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"
import ALSU_sequencer_pkg::*;
import ALSU_sequence_item_pkg::*;

class alsu_main_sequence extends uvm_sequence #(alsu_seq_item);
    `uvm_object_utils(alsu_main_sequence);
    alsu_seq_item item;

    function new(string name = "alsu_main_sequence");
        super.new(name);
    endfunction

    task body;
        repeat(1000) begin
            item = alsu_seq_item::type_id::create("item");
            start_item(item);
            assert(item.randomize());
            finish_item(item);
        end
    endtask
endclass
endpackage